library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity controlMemory is
 	
 	port (
			Input : in std_logic_vector(7 downto 0);

			controlWord : out std_logic_vector(27 downto 0)
		);

 end entity controlMemory; 


architecture Behavioral of controlMemory is
 type mem_array is array(0 to 255) of std_logic_vector(27 downto 0);

 begin
	memory_m: process(Input)
		variable control_mem : mem_array:=(
			-- 0
			x"1020304", --0
            x"1020224", --1
            x"102000C", --2
            x"1020001", --3
            x"1020014", --4
            x"10200E4", --5
            x"1020024", --6
            x"122A002", --7
            x"17E2002", --8
            x"0000000", --9 
            x"0000000", --A 
            x"0000000", --B 
            x"0000000", --C 
            x"0000000", --D 
            x"0000000", --E 
            x"0000000", --F

    		-- 1
            x"110C002", --0
            x"0030000", --1
            x"112A002", --2
            x"0000000", --3 
            x"0000000", --4 
            x"0000000", --5 
            x"0000000", --6 
            x"18FA002", --7
            x"113C002", --8 
            x"0000000", --9 
            x"0000000", --A
            x"0000000", --B 
            x"0000000", --C 
            x"0000000", --D 
            x"0000000", --E 
            x"0000000", --F
 			-- 2
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- 3
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- 4
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- 5
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- 6
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- 7
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- 8
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- 9
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- a
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- b
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- c
			x"C10C002", -- 0
	        x"0030000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- d
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- e
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000", -- F
 			-- f
			X"0000000", -- 0
			X"0000000", -- 1
			X"0000000", -- 2
			X"0000000", -- 3
			X"0000000", -- 4
			X"0000000", -- 5
			X"0000000", -- 6
			X"0000000", -- 7
			X"0000000", -- 8
			X"0000000", -- 9
			X"0000000", -- A
			X"0000000", -- B
			X"0000000", -- C
			X"0000000", -- D
			X"0000000", -- E
			X"0000000" -- F
		);

		variable addr : integer;
	begin	
		addr := conv_integer(Input);
		controlWord <= control_mem(addr);
	end process;	

end Behavioral;

