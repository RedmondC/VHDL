library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity MemoryM is
 	
 	port (
			InputIndex : in std_logic_vector(15 downto 0);
			dataIn : in std_logic_vector(15 downto 0);
			MW : in std_logic;
			dataOut : out std_logic_vector(15 downto 0)
		);

 end entity MemoryM; 


architecture Behavioral of MemoryM is
 type mem_array is array(0 to 511) of std_logic_vector(15 downto 0);

 begin
	memory_m: process(InputIndex,dataIn,MW)
		variable Memory : mem_array:=(
			x"0000", --0 
        x"0000", --1 Reg0 = 0
        x"0041", --2 ...
        x"0082", --3 ...
        x"00C3", --4 ...
        x"0104", --5 ...
        x"0145", --6 ...
        x"0186", --7 ...
        x"01C7", --8 Reg7 = 7
        x"024A", --9 ADI : Reg1 = Reg1 + 2
        x"0410", --A LDR : load 0x41 to Reg0
        x"0601", --B STR : store R1 into memory
        x"09D0", --C INC : Reg7 = Reg2 + 1
        x"0BF8", --D NOT : NOT value in Reg7
        x"0C91", --E ADD : Reg2 = Reg2 + Reg1
        x"0E12", --F B   : Branch past next instruction

        --module 01
        x"0000", --0 Should be skipped
        x"0040", --1 Reg1 = 0
        x"1002", --2 BNZ : branch conditionally if Z is not set
        x"01C7", --3 Should be skipped
        x"0041", --4 R1 = 1
        x"0000", --5 R0 = 0 forever
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 03
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 04
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 05
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 06
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 07
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 08
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 09
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 0a
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 0b
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 0c
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 0d
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
			-- 0e
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 0f
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
			-- 10
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
			-- 11
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 12
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 13
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 14
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 15
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 16
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 17
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 18
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 19
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 1a
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 1b
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 1c
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 1d
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 1e
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", -- F
 			-- 1f
			X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000" -- F
		);

		variable addr : integer range 0 to 511;
		variable addressOut : std_logic_vector(15 downto 0);
	begin	
		addr := conv_integer(InputIndex(8 downto 0));
		addressOut := Memory(addr);

		if MW = '1' then
        	Memory(addr) := dataIn;
        else
			dataOut <= addressOut;
		end if;	
							
		dataOut <= Memory(addr);
	end process;	

 end Behavioral;

